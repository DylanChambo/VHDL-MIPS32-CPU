package types is
    type ALUControl is (ALU_AND, ALU_OR, ALU_ADD, ALU_SUB, ALU_SLT);
end package types;