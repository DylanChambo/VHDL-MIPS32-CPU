library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity write_back is
    port (
        I_CLK : in std_logic;
        I_RST : in std_logic
    );
end write_back;

architecture behavioural of write_back is

begin

end architecture;