library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity register_file is
    port (
        I_CLK : in std_logic;
        I_RST : in std_logic
    );
end register_file;

architecture behavioural of register_file is

begin

end architecture;