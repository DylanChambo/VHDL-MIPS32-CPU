library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity data_mem is
    port (
        I_CLK : in std_logic;
        I_RST : in std_logic
    );
end data_mem;

architecture behavioural of data_mem is

begin

end architecture;