library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.types.all;

entity control is
    port (
        I_CLK : std_logic
    );
end control;

architecture behavioural of control is

begin

end architecture;