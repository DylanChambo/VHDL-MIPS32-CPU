library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity forwarding_unit is
    port (
        I_CLK : in std_logic;
        I_RST : in std_logic
    );
end forwarding_unit;

architecture behavioural of forwarding_unit is

begin

end architecture;