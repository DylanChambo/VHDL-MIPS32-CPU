library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity hazard_detection_unit is
    port (
        I_CLK : in std_logic;
        I_RST : in std_logic
    );
end hazard_detection_unit;

architecture behavioural of hazard_detection_unit is

begin

end architecture;